module template_tb;
//===========================================================================
// REG and WIRE declaration
//===========================================================================
reg clk;
reg rst;


//===========================================================================
// Device Under Test
//===========================================================================
template dut(
  .clk(clk),
  .rst(rst),



);

//===========================================================================
// Always blocks
//===========================================================================
always
  #6.25 clk = !clk;


//===========================================================================
// initial blocks
//===========================================================================
initial begin





end



endmodule
