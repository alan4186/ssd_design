`timescale 1ns/10ps
module crc_buffer_tb;
//===========================================================================
// REG and WIRE declaration
//===========================================================================
reg clk;
reg rst;
reg [7:0] data;
reg rdreq;
reg wrreq;

wire empty;
wire full;
wire [7:0] q;

//===========================================================================
// Device Under Test
//===========================================================================
crc_buffer dut(
  .clock(clk),
  .aclr(!rst),
  .data(data),
  .rdreq(rdreq),
  .wrreq(wrreq),
  .empty(empty),
  .full(full),
  .q(q)

);

//===========================================================================
// Always blocks
//===========================================================================
always
  #5 clk = !clk;


//===========================================================================
// initial blocks
//===========================================================================
initial begin
  clk = 1'b1;
  rst = 1'b1;
  data = 8'd0;
  rdreq = 1'd0;
  wrreq = 1'd0;

  #10
  rst = 1'b0;
  #10
  rst = 1'b1;
  #20
  wrreq = 1'd1;
  #40
  wrreq = 1'd0;

  #100
  $stop;



end



endmodule
